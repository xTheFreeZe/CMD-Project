// V Template
// Run this code with: v run main.v
// Generate the binary by either running: v -prod -o main main.v or v .
module main

fn main() {
	println('Hello, World!')
}
